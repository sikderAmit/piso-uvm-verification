package my_pkg;

//tb-files including
piso_intf.sv
piso_seq_item.sv
piso_sequence.sv

piso_mntr.sv
piso_drvr.sv
piso_predictor.sv
piso_scb.sv
piso_agnt.sv
piso_env.sv

piso_test.sv
tb_top.sv

endpackage